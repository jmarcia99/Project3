`ifndef AES_CORE_H
  `define AES_CORE_H

  `define DRV_CB aes_vif.aes_drv_cb
  `define MON_CB aes_vif.aes_mon_cb
`endif
