/* 
* AES Core to UART Transmitter Testbench
* Created By: Jordi Marcial Cruz
* Project: AES-128 Encryption Core
* Updated: May 17th, 2025
*
* Description:
* This testbench verifies the full data path from AES encryption
* to serial transmission via UART. It connects the AES-128 Core, Output Buffer,
* and UART Transmitter modules through interface-bound signals.
*
* Testbench Highlights:
* - Provides class-based infrastructure for stimulus generation, driving, monitoring,
*   and scoreboarding.
* - Utilizes a software-style reference model to validate the AES encryption against DUT output.
* - Captures UART serial output byte-by-byte, reassembles it, and compares with the
*   encrypted text generated by the reference model.
* - Supports deterministic test cases, randomized vector injection, and stress testing.
*/

`include "AES_Core_Uart.svh"
`timescale 1ns/10ps

import TestbenchPkg::*;

// =============================
// ReferenceModel Class
// Provides model of AES encryption
// =============================
class ReferenceModel extends RefModelPkg::TextEncryption;
  function void f_initial_report();
    $display("Reference model created");
  endfunction

  function new();
    f_initial_report();
  endfunction

  function void f_set_debug();
    this.debug_key_exp = 0;
    $display("---Debug set, showing all expected keys---");
  endfunction

  function void f_encrypt_plain_text (
    input key_t original_key,
    input key_t plain_text
  );
    this.key = original_key;
    this.round_key[0] = original_key;
    this.state_text = plain_text;
    super.f_expand_key(); 
    super.f_encrypt_text();
  endfunction 
endclass : ReferenceModel

// =============================
// Packet Class
// Stores and tracks input stimulus (AES Key and Plaintext)
// =============================
class Packet extends TestbenchPkg::Packet;
  rand pkt_key_t key_pkt;
  rand pkt_text_t text_pkt;

  function void f_create_packet (
    input pkt_key_t key_pkt,
    input pkt_text_t text_pkt
  );
    this.key_pkt = key_pkt;
    this.text_pkt = text_pkt;
    this.pkt_count++;
  endfunction

  function void f_initial_report();
    $display("[%0d][GEN] Packet generated", $stime);
  endfunction

  function void post_randomize();
    this.pkt_count++;
  endfunction
endclass : Packet

// =============================
// Sample Class
// Captures UART byte-level output reconstructed from serial stream
// =============================
class Sample extends TestbenchPkg::Sample;
  logic [7:0] serial_smpl;

  function new (logic [7:0] serial_smpl);
    this.serial_smpl = serial_smpl;
    this.smpl_count++;
    f_initial_report();
  endfunction

  function void f_initial_report();
    if (smpl_count == 16) begin 
      $display("[%0d][MON] All 16 Samples put into Monitor Mailbox", $stime);
      smpl_count = 0;
    end
  endfunction
endclass : Sample

// =============================
// Generator Class
// Randomizes and creates AES key/plaintext packets
// =============================
class Generator extends TestbenchPkg::Generator;
  Packet pkt;

  function new(mailbox generator_mbx);
    this.generator_mbx = generator_mbx;
    f_initial_report();
  endfunction

  function void f_initial_report();
    $display("Generator instantiated in testbench");
  endfunction

  task t_generate_pkts(input int num_of_pkts);
    $display("[%0d] Generating %0d randomized packets", $stime, num_of_pkts);
    repeat (num_of_pkts) begin
      pkt = new();
      pkt.randomize();
      generator_mbx.put(pkt);
    end
    $display("[%0d] %0d Packets put into Generator Mailbox", $stime, num_of_pkts);
  endtask

  task t_create_pkt (
    input pkt_key_t key,
    input pkt_text_t text
  );
    $display("[%0d][GEN] Creating packet", $stime);
    pkt = new();
    pkt.f_create_packet(key, text);
    generator_mbx.put(pkt);
    $display("[%0d][GEN] Packet put into Generator Mailbox", $stime);
  endtask
endclass : Generator

// =============================
// Scoreboard Class
// Assembles and validates received UART data against AES reference
// =============================
class Scoreboard extends TestbenchPkg::Scoreboard;
  ReferenceModel ref_model;
  smpl_text_t expected_text;
  Packet pkt;
  Sample smpl;
  static int pkts_read;

  logic [0:15][7:0] assembled_smpl;
  int smpl_index;

  function new (
    ReferenceModel ref_model,
    mailbox driver_mbx,
    mailbox monitor_mbx
  );
    this.ref_model = ref_model;
    this.driver_mbx = driver_mbx;
    this.monitor_mbx = monitor_mbx;
    this.smpl_index = 0;
    this.errors = 0;
    this.pkts_read = 0;
    f_initial_report();
  endfunction

  function void f_initial_report(); 
    $display("Scoreboard instantiated in testbench");
  endfunction

  task t_run();
    forever begin
      driver_mbx.get(pkt);

      repeat(16) begin
        monitor_mbx.get(smpl);
        assembled_smpl[smpl_index] = smpl.serial_smpl;
        smpl_index++;
      end

      t_check_results(); 
    end
  endtask

  task t_check_results();
    expected_text = f_retreive_expected_text(pkt.key_pkt, pkt.text_pkt);

    if (expected_text !== assembled_smpl) begin
      $display("[%0d][SB] Expected Text: %h, Received Text: %h", $stime, expected_text, assembled_smpl);
      errors++;
    end else begin
      $display("[%0d][SB] Text Received: %h", $stime, assembled_smpl);
      $display("[%0d][SB] Text Expected: %h \n", $stime, expected_text);
    end

    pkts_read++;
    smpl_index = 0;
    assembled_smpl = 0;
  endtask

  function pkt_text_t f_retreive_expected_text (
    input pkt_key_t key,
    input pkt_text_t text
  );
    ref_model.f_encrypt_plain_text(key, text);
    return ref_model.state_text;
  endfunction

  function void f_final_report();
    if (errors > 0) 
      $display("[SB] Testbench FAILED with %0d errors!", errors);
    else if (pkts_read !== pkt.pkt_count) 
      $display("[SB] Testbench FAILED all packets not received!");
    else
      $display("[SB] Testbench PASSED with 0 errors! Received all %0d packets!", pkts_read); 
  endfunction
endclass : Scoreboard

// =============================
// Driver Class
// Drives encryption inputs into AES Core
// =============================
class Driver extends TestbenchPkg::Driver;
  virtual AES_Core_Interface.AES_Driver aes_vif;
  Packet pkt;
  int debug;

  function new (
    virtual AES_Core_Interface.AES_Driver aes_vif,
    mailbox driver_mbx,
    mailbox generator_mbx
  );
    this.aes_vif = aes_vif;
    this.driver_mbx = driver_mbx;
    this.generator_mbx = generator_mbx;
    this.debug = 0;
  endfunction

  function void f_initial_report();
    $display("Driver instantiated in testbench");
  endfunction

  task t_initialize_signals();
    `DRV_CB.start_encryption <= 0;
    `DRV_CB.plain_text <= 0;
    `DRV_CB.original_key <= 0;
  endtask

  task t_run();
    forever begin
      @(`DRV_CB);
      if (!`DRV_CB.output_buffer_full) begin 
        generator_mbx.get(pkt);
        driver_mbx.put(pkt);
        `DRV_CB.start_encryption <= 1;
        `DRV_CB.plain_text <= pkt.text_pkt;
        `DRV_CB.original_key <= pkt.key_pkt;
        if (debug) $display("[%0d][DRV] Sending -> Key: %h, Plain Text: %h", $stime, pkt.key_pkt, pkt.text_pkt);
        else       $display("[%0d][DRV] Text Packet Sent", $stime);
        @(`DRV_CB);
        `DRV_CB.start_encryption <= 0;
        `DRV_CB.plain_text <= 0;
        `DRV_CB.original_key <= 0;
        repeat(11) @(`DRV_CB);
      end
    end
  endtask
endclass : Driver

// =============================
// Monitor Class
// Shifts out received UART bytes and sends to scoreboard
// =============================
class Monitor extends TestbenchPkg::Monitor;
  virtual Uart_Interface.Tx_Monitor uart_vif;
  const int CLKS_PER_BIT;
  Sample smpl;

  logic [7:0] return_shift_register;
  int debug;

  function new (
    virtual Uart_Interface.Tx_Monitor uart_vif,
    int CLKS_PER_BIT,
    mailbox monitor_mbx
  );
    this.uart_vif = uart_vif;
    this.monitor_mbx = monitor_mbx;
    this.return_shift_register = '0;
    this.CLKS_PER_BIT = CLKS_PER_BIT;
    this.debug = 0;
    f_initial_report();
  endfunction 

  function void f_initial_report(); 
    $display("Monitor instantiated in testbench");
  endfunction

  task t_run();
    forever begin 
      if (`MON_CB.tx_active) begin 
        @(`MON_CB);

        fork 
          begin 
            repeat(CLKS_PER_BIT) @(`MON_CB);

            repeat(8) begin 
              return_shift_register[7:0] <= {`MON_CB.tx_serial_out, return_shift_register[7:1]};
              repeat(CLKS_PER_BIT) @(`MON_CB); 
            end 

            return_shift_register <= return_shift_register;
            @(`MON_CB);

            if (debug) $display("[%0d][MON] Received -> Serial Data: %h", $stime, return_shift_register);

            smpl = new(return_shift_register);
            monitor_mbx.put(smpl);
          end

          begin 
            while (!`MON_CB.tx_done) @(`MON_CB);
          end
        join

      end else begin 
        @(`MON_CB);
      end
    end
  endtask
endclass : Monitor

  
// ============================= 
// Testbench Top Level 
// =============================
module AES_Core_to_Uart_TB ();
  
  localparam CLOCK_PERIOD = 500; // 50 MHz clock
  localparam CLKS_PER_BIT = 434; // 50000000 / 115200 = 434 Clocks Per Bit.
  localparam DATA_WIDTH = 128;   // AES Block Size
   
  logic clk;
  logic reset_n;
  
  logic start_encrypt;
  text_t provided_text;
  key_t provided_key;
  
  logic uart_serial_out;
  logic uart_buffer_full;
  logic text_ready;
  text_t cipher_text;
  
  AES_Core_Interface aes_if (
    .clk				(clk),
    .reset_n			(reset_n),
    .start_encrypt		(start_encrypt),
    .output_buffer_full	(uart_buffer_full),
    .provided_text		(provided_text),
    .provided_key		(provided_key),
    .final_text			(cipher_text),
    .finished_encrypt	(text_ready)
  );
  
  Key_Expansion Key_Exp (
    .kx_if			(aes_if)
  );
  
  SBox SBox_Tables (
    .sb_if			(aes_if)
  );
  
  Shift_Rows Shift_Rows (
    .sr_if			(aes_if) 
  );
  
  Mix_Columns Mix_Columns (
    .mc_if			(aes_if)
  );
  
  AES_Controller Controller (
    .cntrl_if		(aes_if)
  );
  
  
  Uart_Interface uart_if (
    .clk				(clk),
    .reset_n			(reset_n),
    .uart_serial_out	(uart_serial_out),
    .uart_buffer_full	(uart_buffer_full),
    .text_ready			(text_ready),
    .cipher_text		(cipher_text)
  );
   
  Uart_Tx #(
    .CLKS_PER_BIT		(CLKS_PER_BIT)
  ) Transmitter (
    .tx_if				(uart_if)
  );
  
  Output_Buffer #(
    .DATA_WIDTH 		(DATA_WIDTH)
  ) Buffer (
    .buff_if			(uart_if)
  );
  
  mailbox generator_mbx;
  mailbox driver_mbx;
  mailbox monitor_mbx;
  ReferenceModel ref_model;
  Generator gen;
  Scoreboard sb;
  Driver drv;
  Monitor mon;

  task t_reset_dut();
    reset_n = 0;
    drv.t_initialize_signals();
    #5;
    reset_n = 1;
  endtask
  
  task t_set_debug(input bit flag); 
    drv.debug = flag;
    mon.debug = flag;
  endtask

  task t_run_processes();
    fork
      drv.t_run();
      mon.t_run();
      sb.t_run();
    join_none
  endtask

  task t_timeout(input int cycles);
    repeat(cycles * CLKS_PER_BIT) @(posedge clk);
    $fatal("Testbench timed out");
  endtask

  task t_send_key_and_text (
    input key_t key,
  	input text_t text
  );
    gen.t_create_pkt(key, text);
  endtask

  task t_send_randomized_pkts(input int num_of_pkts);
    gen.t_generate_pkts(num_of_pkts);
  endtask
  
  default clocking cb @(posedge clk); endclocking
 
  initial begin 
    clk = 1;
    forever #(CLOCK_PERIOD/2) clk = ~clk;
  end
   
  // Main Testing:
  initial begin 
    ref_model = new;
    driver_mbx = new; 
    monitor_mbx = new;
    generator_mbx = new; 
    gen = new(generator_mbx);
    sb = new(ref_model, driver_mbx, monitor_mbx);
    drv = new(aes_if, driver_mbx, generator_mbx);
    mon = new(uart_if, CLKS_PER_BIT, monitor_mbx);
    
    $display("Beginning testbench, initializing signals...");
    t_reset_dut();
    t_set_debug(1);

    fork
      t_timeout(55000);
      t_run_processes();
    join_none

    // Test vectors from CSRC
    $display("Beginning Direct Test Cases...");
    t_send_key_and_text(128'h000102030405060708090a0b0c0d0e0f, 128'h00112233445566778899aabbccddeeff);
    t_send_key_and_text(128'h139a35422f1d61de3c91787fe0507afd, 128'hb9145a768b7dc489a096b546f43b231f);
    t_send_key_and_text(128'hc459caeebf2c42586c01666a9334b97b, 128'hd7c3ffac9031238650901e157364c386);
    t_send_key_and_text(128'h786ffd349283cd971069dd42527719df, 128'hbc3637da2daf8fcf7c68bb28c143a0a4);
    t_send_key_and_text(128'he4e755efeb0c85480aad4e28a8e28773, 128'h9c88a8db798f48df1ac4936afa959eac);
    t_send_key_and_text(128'h2573ded4a95abd8ab3250cecebc5bb29, 128'h79ee212734f14d1bf5a59d46e8c2fa34);
    t_send_key_and_text(128'he98ef4285586a1b458427105b4712e42, 128'hc52263efa6379209d17e87ac250615cb);
    t_send_key_and_text(128'hdae519292b9603f3b6d0e99dd6323f21, 128'h336bed017e10a247ee92989862431163);
    t_send_key_and_text(128'h6bd60971346858e31c3f37254f18d339, 128'hb13310581ffe5b10aaefdeb8992aec18);
    t_send_key_and_text(128'hdb3ce492c786e70c94bd1d4b91018388, 128'hb0eaede3f3eebfef88822a6ede1950b1);
    
    $display("\nBeginning Random Test Cases...");
    t_send_randomized_pkts(30);
    
    repeat (3500) ##CLKS_PER_BIT;
    
    $display("\nBeginning Stress Test, bombarding output buffer...");
    t_set_debug(0);
    t_send_randomized_pkts(250);

    repeat (50000) ##CLKS_PER_BIT;
    sb.f_final_report();
    $finish;  
    
    end
endmodule























































 










