`ifndef KEY_EXPANSION_H
  `define KEY_EXPANSION_H

  `define DRV_CB aes_vif.kx_drv_cb
  `define MON_CB aes_vif.kx_mon_cb
`endif
