`ifndef UART_TX_H
  `define UART_TX_H

  `define DRV_CB uart_vif.tx_drv_cb
  `define MON_CB uart_vif.tx_mon_cb
`endif
