`ifndef AES_CORE_UART_H
  `define BUFFERED_UART_H

  `define DRV_CB aes_vif.aes_drv_cb
  `define MON_CB uart_vif.tx_mon_cb
`endif
